module alu_4bit
  (input sel,
   input left_operand,
   input right_operand,
   output result
